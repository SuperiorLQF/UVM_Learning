module MCHDP(
	input 	clk,
	input	rst_n,
	input	[7:0]	sop,
	input	[7:0]	eop,
	input	[7:0]	vld,
	input	[95:0]	in_chan_data
);
endmodule